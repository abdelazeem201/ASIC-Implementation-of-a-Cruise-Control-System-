* Nettran: AMD.64 Release B-2008.09.SP5.26004 2012/07/19
* Created:  12/20/2017   8:49
* Options: -rootCell cruisecontrol -verilog-b0 VSS -verilog-b1 VDD -sp /home/standard_cell_libraries/NangateOpenCellLibrary_PDKv1_3_v2010_12/lib/Back_End/spice/NangateOpenCellLibrary.spi -verilog ../../../pnr/output/cruisecontrol_icc.v -outType spice -outName cruisecontrl.sp 

.GLOBAL VDD VSS 

.SUBCKT TAP VDD VSS 
.ENDS

.SUBCKT XOR2_X2 A B Z VDD VSS 
M_i_41_29 net_003 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_47_27 Z A net_003 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_53_18 net_003 B Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_53 net_003 B Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_47 Z A net_003 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_41 net_003 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_35 VDD B net_002 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_30 net_002 A net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_35 Z net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_19_23 net_001b A Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_24_4 VSS B net_001b VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_24 VSS B net_001 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_19 net_001 A Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_13 Z net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 VSS B net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_000 A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT XNOR2_X2 A B ZN VDD VSS 
M_i_53 VDD B net_003 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_53_25 VDD B net_003b VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_48_8 net_003b A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_48 net_003 A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_29 net_000 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_36 VDD B net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_42 ZN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_42_14 ZN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_23 net_002 B ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_23_12 net_002 B ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_17 ZN A net_002 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_17_20 ZN A net_002 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_001 A net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS B net_001 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_11 net_002 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_11_23 net_002 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT TLAT_X1 D G OE Q VDD VSS 
M_i_111 Q net_005 net_010 VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_106 net_010 net_003 VDD VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_91 net_005 OE VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_99 VDD net_003 net_006 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_85 VDD net_006 net_009 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_81 net_009 net_001 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_75 net_003 net_000 net_008 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_70 net_008 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_64 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_57 VDD G net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_51 Q OE net_007 VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_47 net_007 net_003 VSS VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_34 net_005 OE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 VSS net_003 net_006 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 VSS net_006 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_000 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_001 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS G net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT TINV_X1 EN I ZN VDD VSS 
M_i_29 ZN EN net_002 VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24 net_002 I VDD VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VDD EN net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_11 ZN net_000 net_001 VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_7 net_001 I VSS VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0 VSS EN net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT TBUF_X8 A EN Z VDD VSS 
M_i_42 VDD EN NEN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1 dummy0 EN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0 x A dummy0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_130 x A dummy0a VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_114 dummy0a EN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_48_94 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64_92 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_48 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_9 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_18 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8_39 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19_50 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VSS EN NEN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_129 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_113 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_47_77 VSS NEN dummy1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63_69 dummy1 A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63 dummy1a A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_47 VSS NEN dummy1a VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_42 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_37 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13_45 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6_40 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
.ENDS

.SUBCKT TBUF_X4 A EN Z VDD VSS 
M_i_42 VDD EN NEN VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_1 dummy0 EN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0 x A dummy0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_48 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VSS EN NEN VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_14 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63 dummy1 A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_47 VSS NEN dummy1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
.ENDS

.SUBCKT TBUF_X2 A EN Z VDD VSS 
M_i_42 VDD EN NEN VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_1_48 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0 VDD A dummy0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1 dummy0 EN x VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VSS EN NEN VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_14_47 VSS NEN dummy1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63 dummy1 A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
.ENDS

.SUBCKT TBUF_X16 A EN Z VDD VSS 
M_i_42 VDD EN NEN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1 dummy0 EN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0 x A dummy0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_130 x A dummy0a VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_114 dummy0a EN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_48_94 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64_92 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_0_64 VDD A y VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24_1_48 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_24 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_9 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_18 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8_39 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19_50 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_10 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_83 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8_42 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19_51 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_9_17 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_18_103 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_8_39_66 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_24_3_19_50_12 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VSS EN NEN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_129 VSS A x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_113 VSS EN x VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_47_77 VSS NEN dummy1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63_69 dummy1 A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15_63 dummy1a A y VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14_47 VSS NEN dummy1a VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_42 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_37 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13_45 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6_40 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_116 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_106 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13_120 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6_43 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_42_108 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_37_112 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_13_45_122 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
M_i_0_6_6_40_125 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
.ENDS

.SUBCKT TBUF_X1 A EN Z VDD VSS 
M_i_42 VDD EN NEN VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_1 dummy0 EN x VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_0 VDD A dummy0 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_1_48 y NEN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24_0_64 VDD A y VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24 VDD y Z VDD PMOS_VTL L=0.050000U W=0.540000U 
M_i_17 VSS EN NEN VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_14 VSS EN x VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_15 VSS A x VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_14_47 VSS NEN dummy1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_15_63 dummy1 A y VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS x Z VSS NMOS_VTL L=0.050000U W=0.355000U 
.ENDS

.SUBCKT SDFF_X2 D SE SI CK Q QN VDD VSS 
M_i_210 net_013 SE VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_204 VDD D net_019 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_200 net_019 SE net_011 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_194 net_011 net_013 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_189 net_018 SI VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_155 VDD net_007 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_176 VDD net_011 net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_172 net_017 net_004 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_166 net_007 net_009 net_016 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_162 net_016 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_182 net_009 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_149 net_004 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 VDD net_007 net_015 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_138 net_015 net_009 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_132 net_002 net_004 net_014 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_128 net_014 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_115_2 QN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_115 QN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_108 VDD net_002 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_108_51 VDD net_002 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_121 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_102 net_013 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_81 net_010 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_86 net_011 net_013 net_010 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_92 net_012 SE net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_96 VSS SI net_012 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_47 VSS net_007 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_69 VSS net_011 net_008 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_64 net_008 net_009 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_58 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_54 net_006 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_75 net_009 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_004 net_009 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_34 VSS net_007 net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_30 net_003 net_004 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_24 net_002 net_009 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_20 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_7_4 QN net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 QN net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS net_002 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_50 VSS net_002 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_13 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT SDFF_X1 D SE SI CK Q QN VDD VSS 
M_i_210 net_013 SE VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_204 VDD D net_019 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_200 net_019 SE net_011 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_194 net_011 net_013 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_189 net_018 SI VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_155 VDD net_007 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_176 VDD net_011 net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_172 net_017 net_004 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_166 net_007 net_009 net_016 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_162 net_016 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_182 net_009 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_149 net_004 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 VDD net_007 net_015 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_138 net_015 net_009 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_132 net_002 net_004 net_014 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_128 net_014 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_121 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_108 VDD net_002 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_115 QN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_102 net_013 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_81 net_010 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_86 net_011 net_013 net_010 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_92 net_012 SE net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_96 VSS SI net_012 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_47 VSS net_007 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_69 VSS net_011 net_008 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_64 net_008 net_009 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_58 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_54 net_006 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_75 net_009 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_004 net_009 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_34 VSS net_007 net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_30 net_003 net_004 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_24 net_002 net_009 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_20 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_13 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS net_002 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 QN net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT SDFFS_X2 D SE SI SN CK Q QN VDD VSS 
M_i_230_17 VDD net_015 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_230 VDD net_015 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_237 Q net_012 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_237_1 Q net_012 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_224 VDD net_012 net_015 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_218 net_015 SN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_189 VDD net_007 net_010 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_212 VDD net_015 net_022 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_208 net_022 net_005 net_012 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_201 net_012 net_004 net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_197 net_021 net_007 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_178 net_019 SN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_172 VDD net_010 net_019 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_168 net_019 net_004 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_162 net_007 net_005 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_157 net_018 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_150 net_005 net_004 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 VDD CK net_004 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_137 VDD SI net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_133 net_017 net_000 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_127 net_002 SE net_016 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_123 net_016 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_116 VDD SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_103_26 VSS net_015 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_103 VSS net_015 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_110 Q net_012 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_110_2 Q net_012 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_97 VSS net_012 net_014 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_93 net_014 SN net_015 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_66 net_010 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_87 VSS net_015 net_013 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_83 net_013 net_004 net_012 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_77 net_012 net_005 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_73 net_011 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_60 VSS SN net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_51 net_008 net_005 net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_45 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_006 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_34 net_005 net_004 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 VSS CK net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 SI VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_11 net_002 SE net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_17 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_21 VSS D net_003 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_0 VSS SE net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT SDFFS_X1 D SE SI SN CK Q QN VDD VSS 
M_i_230 VDD net_015 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_237 Q net_012 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_224 VDD net_012 net_015 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_218 net_015 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_212 VDD net_015 net_022 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_208 net_022 net_005 net_012 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_201 net_012 net_004 net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_197 net_021 net_007 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_189 VDD net_007 net_010 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_178 net_019 SN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_172 VDD net_010 net_019 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_168 net_019 net_004 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_162 net_007 net_005 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_157 net_018 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_150 net_005 net_004 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 VDD CK net_004 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_137 VDD SI net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_133 net_017 net_000 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_127 net_002 SE net_016 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_123 net_016 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_116 VDD SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_103 VSS net_015 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_110 Q net_012 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_97 net_015 net_012 net_014 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_93 net_014 SN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_87 VSS net_015 net_013 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_83 net_013 net_004 net_012 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_77 net_012 net_005 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_73 net_011 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_66 net_010 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_60 VSS SN net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_51 net_008 net_005 net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_45 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_006 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_34 net_005 net_004 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 VSS CK net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 SI VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_11 net_002 SE net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_17 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_21 VSS D net_003 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_0 VSS SE net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT SDFFR_X2 D RN SE SI CK Q QN VDD VSS 
M_i_236 net_015 SE VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_230 VDD D net_022 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_226 net_022 SE net_013 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_220 net_013 net_015 net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_215 net_021 SI VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_181 VDD RN net_006 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_174 net_006 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_203 VDD net_013 net_020 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_199 net_020 net_005 net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_193 net_009 net_011 net_019 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_188 net_019 net_006 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_167 VDD net_011 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_209 net_011 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_157 net_018 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_161 net_003 net_011 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_146 net_017 net_005 net_003 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_151 VDD net_000 net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_136 net_017 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_116_1 VDD net_000 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_116 VDD net_000 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_123 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_123_146 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_129 VDD net_003 net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_110 net_015 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_89 net_012 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_94 net_013 net_015 net_012 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_100 net_014 SE net_013 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_104 VSS SI net_014 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_56 VSS RN net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_51 net_007 net_009 net_006 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_77 VSS net_013 net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_72 net_010 net_011 net_009 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_66 net_009 net_005 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_62 net_008 net_006 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_45 net_005 net_011 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_83 net_011 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_39 VSS net_009 net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_35 net_004 net_005 net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_29 net_003 net_011 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_25 net_002 net_000 net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_21 net_001 RN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_10 VSS net_000 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS net_000 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7_145 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_13 VSS net_003 net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT SDFFR_X1 D RN SE SI CK Q QN VDD VSS 
M_i_236 net_015 SE VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_230 VDD D net_022 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_226 net_022 SE net_013 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_220 net_013 net_015 net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_215 net_021 SI VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_181 VDD RN net_006 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_174 net_006 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_203 VDD net_013 net_020 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_199 net_020 net_005 net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_193 net_009 net_011 net_019 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_188 net_019 net_006 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_167 VDD net_011 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_209 net_011 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_157 net_018 net_009 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_161 net_003 net_011 net_018 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_146 net_017 net_005 net_003 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_151 VDD net_000 net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_136 net_017 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_129 VDD net_003 net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_123 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_116 VDD net_000 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_110 net_015 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_89 net_012 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_94 net_013 net_015 net_012 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_100 net_014 SE net_013 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_104 VSS SI net_014 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_56 VSS RN net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_51 net_007 net_009 net_006 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_77 VSS net_013 net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_72 net_010 net_011 net_009 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_66 net_009 net_005 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_62 net_008 net_006 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_45 net_005 net_011 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_83 net_011 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_39 VSS net_009 net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_35 net_004 net_005 net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_29 net_003 net_011 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_25 net_002 net_000 net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_21 net_001 RN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_13 VSS net_003 net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS net_000 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT SDFFRS_X2 D RN SE SI SN CK Q QN VDD VSS 
M_i_138 VDD SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_145 net_020 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_149 net_002 SE net_020 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_155 net_021 net_000 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_159 VDD SI net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_183 VDD net_002 net_022 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_178 net_022 net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_193 net_007 net_004 net_023 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_189 net_023 net_010 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_203 VDD SN net_023 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_172 net_005 net_004 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_211 net_010 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_217 VDD net_007 net_010 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_228 VDD net_007 net_025 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_223 net_025 net_004 net_013 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_238 net_013 net_005 net_026 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_234 net_026 net_017 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_248 VDD RN net_026 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_165 VDD CK net_004 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_262 VDD net_013 net_017 VDD PMOS_VTL L=0.050000U W=0.485000U 
M_i_255 net_017 SN VDD VDD PMOS_VTL L=0.050000U W=0.485000U 
M_i_270 net_019 RN VDD VDD PMOS_VTL L=0.050000U W=0.485000U 
M_i_284 VDD net_017 net_019 VDD PMOS_VTL L=0.050000U W=0.485000U 
M_i_277_67 VDD net_017 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_277 VDD net_017 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_290 Q net_019 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_290_11 Q net_019 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 VSS SE net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_22 VSS D net_003 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_12 net_002 SE net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 SI VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_41 net_006 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_46 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_52 net_008 net_005 net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_60 VSS SN net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_35 net_005 net_004 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_66 net_011 RN net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_71 VSS net_007 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_77 net_012 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_81 net_013 net_005 net_012 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_87 net_014 net_004 net_013 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_015 net_017 net_014 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_95 VSS RN net_015 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 VSS CK net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_101 net_016 net_013 VSS VSS NMOS_VTL L=0.050000U W=0.310000U 
M_i_106 net_017 SN net_016 VSS NMOS_VTL L=0.050000U W=0.310000U 
M_i_119 net_019 RN net_018 VSS NMOS_VTL L=0.050000U W=0.310000U 
M_i_114 net_018 net_017 VSS VSS NMOS_VTL L=0.050000U W=0.310000U 
M_i_125_68 VSS net_017 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_125 VSS net_017 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_132 Q net_019 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_132_2 Q net_019 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT SDFFRS_X1 D RN SE SI SN CK Q QN VDD VSS 
M_i_138 VDD SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_145 net_020 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_149 net_002 SE net_020 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_155 net_021 net_000 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_159 VDD SI net_021 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_183 VDD net_002 net_022 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_178 net_022 net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_193 net_007 net_004 net_023 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_189 net_023 net_010 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_203 VDD SN net_023 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_172 net_005 net_004 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_211 net_010 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_217 VDD net_007 net_010 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_228 VDD net_007 net_025 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_223 net_025 net_004 net_013 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_238 net_013 net_005 net_026 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_234 net_026 net_017 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_248 VDD RN net_026 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_165 VDD CK net_004 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_262 VDD net_013 net_017 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_255 net_017 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_270 net_019 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_284 VDD net_017 net_019 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_277 VDD net_017 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_290 Q net_019 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 VSS SE net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_22 VSS D net_003 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_12 net_002 SE net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 SI VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_41 net_006 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_46 net_007 net_004 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_52 net_008 net_005 net_007 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_56 net_009 net_010 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_60 VSS SN net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_35 net_005 net_004 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_66 net_011 RN net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_71 VSS net_007 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_77 net_012 net_007 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_81 net_013 net_005 net_012 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_87 net_014 net_004 net_013 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_015 net_017 net_014 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_95 VSS RN net_015 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 VSS CK net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_106 net_017 net_013 net_016 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_101 net_016 SN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_114 net_018 RN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_119 net_019 net_017 net_018 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_125 VSS net_017 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_132 Q net_019 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR4_X4 A1 A2 A3 A4 ZN VDD VSS 
M_i_1_3 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 VDD A4 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 net_2__m1 A3 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 net_1__m1 A2 net_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_0__m1 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN_neg A1 net_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 net_0__m0_0 A2 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 net_1__m0_0 A3 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 net_2__m0_0 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_3 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m1 VSS A4 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 ZN_neg A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 VSS A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 ZN_neg A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 VSS A3 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m0 ZN_neg A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR4_X2 A1 A2 A3 A4 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD A4 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_2 A3 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_1 A2 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS A4 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 ZN_neg A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR3_X4 A1 A2 A3 ZN VDD VSS 
M_i_1_3 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 VDD A3 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_1__m1 A2 net_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 net_0__m1 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN_neg A1 net_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_0__m0_0 A2 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 net_1__m0_0 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_3 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 VSS A3 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 ZN_neg A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 VSS A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 ZN_neg A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR3_X2 A1 A2 A3 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A3 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_1 A2 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS A3 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 ZN_neg A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR2_X4 A1 A2 ZN VDD VSS 
M_i_1_0_x4_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_3 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_2 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_m2__m0 VDD A2 net_0__m0_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_m2__m0 net_0__m0_0__m0_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_m2__m1 ZN_neg A1 net_0__m0_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_m2__m1 net_0__m0_0__m1 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x4_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_3 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_2 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_x2__m0 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_x2__m0 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_x2__m1 VSS A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_x2__m1 ZN_neg A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR2_X2 A1 A2 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 VDD A2 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI33_X1 A1 A2 A3 B1 B2 B3 ZN VDD VSS 
M_i_8 VDD A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 ZN B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 net_3 B2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11 net_4 B3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2 ZN A3 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_0 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 net_0 B3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI22_X4 A1 A2 B1 B2 ZN VDD VSS 
M_i_5__m3 VDD A2 net_1__m3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m3 net_1__m3 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 ZN A1 net_1__m2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m2 net_1__m2 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 VDD A2 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_1__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN A1 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 net_1__m0_0 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m3 VDD B2 net_2__m3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m3 net_2__m3 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m2 ZN B1 net_2__m2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m2 net_2__m2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 VDD B2 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_2__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN B1 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 net_2__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m3 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 ZN A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m3 net_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m3 VSS B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m2 net_0 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m2 VSS B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 VSS B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_0 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI22_X2 A1 A2 B1 B2 ZN VDD VSS 
M_i_5__m1 VDD A2 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_1__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN A1 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 net_1__m0_0 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 VDD B2 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_2__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN B1 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 net_2__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 VSS B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_0 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI222_X4 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_15_3_x4_1 VDD ZN_6 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_0 ZN ZN_6 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_2 VDD ZN_6 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_3 ZN ZN_6 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x2_1 VDD ZN_5 ZN_6 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x2_0 ZN_6 ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11 VDD C2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 net_4 C1 ZN_5 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 ZN_5 B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 net_3 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 A1 ZN_5 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_14_0_x4_3 VSS ZN_6 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_1 ZN ZN_6 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_2 VSS ZN_6 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_0 ZN ZN_6 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_1_x2_0 VSS ZN_5 ZN_6 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_1_x2_1 ZN_6 ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS C2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 net_1 C1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 ZN_5 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN_5 A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI222_X2 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_6__m1 ZN A1 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 net_2__m1 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD A2 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_2__m0_0 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 ZN B1 net_3__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 net_3__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 VDD B2 net_3__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 net_3__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10__m0 ZN C1 net_4__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11__m0 net_4__m0_0 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11__m1 VDD C2 net_4__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10__m1 net_4__m1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0__m1 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1 B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_0 B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_1 B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_0 B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 net_1 C1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m0 VSS C2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m1 net_1 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 VSS C1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI222_X1 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_6 ZN A1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_3 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 ZN C1 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11 net_4 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_0 B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS C1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 net_1 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI221_X4 A B1 B2 C1 C2 ZN VDD VSS 
M_i_13_3_x4_0 VDD ZN_5 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_3_x4_1 ZN ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_3_x4_2 VDD ZN_5 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_3_x4_3 ZN ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_1_x2_0 VDD ZN_4 ZN_5 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_1_x2_1 ZN_5 ZN_4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_3 B1 ZN_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 ZN_4 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 VDD C2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_2 C1 ZN_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_12_0_x4_3 VSS ZN_5 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_2 ZN ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_1 VSS ZN_5 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_0 ZN ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_0_x2_1 VSS ZN_4 ZN_5 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_0_x2_0 ZN_5 ZN_4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 C2 ZN_4 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN_4 C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI221_X2 A B1 B2 C1 C2 ZN VDD VSS 
M_i_7_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 ZN B1 net_3__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 net_3__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 VDD B2 net_3__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 net_3__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 VDD C2 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 net_2__m1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN C1 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_2__m0_0 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_0 net_0 A net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_1 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 VSS B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 net_1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 net_1 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_0 C2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI221_X1 A B1 B2 C1 C2 ZN VDD VSS 
M_i_5 ZN C1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 ZN B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 net_3 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 A net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI21_X4 A B1 B2 ZN VDD VSS 
M_i_4__m3 VDD B2 net_1__m3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m3 net_1__m3 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m2 ZN B1 net_1__m2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 net_1__m2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 VDD B2 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 net_1__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0 ZN B1 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 net_1__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m3 net_0 B2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 ZN B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 net_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 ZN B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_0 B2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_3 net_0 A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_2 VSS A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 net_0 A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 VSS A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI21_X2 A B1 B2 ZN VDD VSS 
M_i_4__m1 VDD B2 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 net_1__m1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0 ZN B1 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 net_1__m0_0 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 net_0 B2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 net_0 A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 VSS A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI211_X4 A B C1 C2 ZN VDD VSS 
M_i_5__m3 VDD C2 net_2__m3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m3 net_2__m3 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 ZN C1 net_2__m2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m2 net_2__m2 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 VDD C2 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_2__m1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN C1 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 net_2__m0_0 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m3 ZN B VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m2 VDD B ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 ZN B VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD B ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m3 net_0 C2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_0 C2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m3 net_0 A net_1__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m3 net_1__m3 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m2 VSS B net_1__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m2 net_1__m2 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_0 A net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_1__m1 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1__m0_0 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI211_X2 A B C1 C2 ZN VDD VSS 
M_i_5__m1 VDD C2 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_2__m1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN C1 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 net_2__m0_0 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 ZN B VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD B ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 net_0 C2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_0 A net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_1__m1 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1__m0_0 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR4_X4 A1 A2 A3 A4 ZN VDD VSS 
M_i_7_1_96 net_2 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_102 net_2 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_1 net_2 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_34_44 net_1 A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_56 net_1 A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_34 net_1 A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_1 A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_88 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_24_95 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_24 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_68 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_6_75 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_6 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_8_108 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3_109 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3_8 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_29_45 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_52 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_29 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_79 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_13_89 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_13 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_77 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_22_71 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_22 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR4_X2 A1 A2 A3 A4 ZN VDD VSS 
M_i_7__m1 VDD A4 net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_2__m1 A3 net_1__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 net_1__m1 A2 net_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_0__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN A1 net_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 net_0__m0_0 A2 net_1__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_1__m0_0 A3 net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 net_2__m0_0 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 VSS A4 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR4_X1 A1 A2 A3 A4 ZN VDD VSS 
M_i_4 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_1 A3 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 ZN A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR3_X4 A1 A2 A3 ZN VDD VSS 
M_i_5_83 net_1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_65 net_1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_56 net_1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_52 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_43 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_34 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_6 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_15 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_24 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_85 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_67 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_58 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_49 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_40 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_31 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_10 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_19 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_28 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR3_X2 A1 A2 A3 ZN VDD VSS 
M_i_5_1_m2__m1 VDD A3 net_1_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_0_m2__m1 net_1_0__m1 A2 net_0_0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1_m2__m1 net_0_0__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1_m2__m0 ZN A1 net_0_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_0_m2__m0 net_0_0__m0_0 A2 net_1_0__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_1_m2__m0 net_1_0__m0_0 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_0_x2__m1 VSS A3 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_1_x2__m1 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x2__m1 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x2__m0 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_1_x2__m0 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0_x2__m0 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR2_X2 A1 A2 ZN VDD VSS 
M_i_3__m0_m2__m1 VDD A2 net_0__m0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m1 net_0__m0__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m0 ZN A1 net_0__m0__m0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_m2__m0 net_0__m0__m0 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m0_x2__m1 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m1 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_x2__m0 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND4_X4 A1 A2 A3 A4 ZN VDD VSS 
M_i_7 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_1 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_52 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_154 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_49 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_100 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6_202 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_87 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_36 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_189 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_15 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_66 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4_168 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 net_2 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3_17 net_2 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3_68 net_2 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3_170 net_2 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 A3 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_43 net_1 A3 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_94 net_1 A3 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_196 net_1 A3 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_75 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_24 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_177 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_34 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_85 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_187 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND4_X2 A1 A2 A3 A4 ZN VDD VSS 
M_i_7__m1 VDD A4 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 ZN A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 VSS A4 net_2__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_2__m1 A3 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_1__m1 A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 A2 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1__m0_0 A3 net_2__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_2__m0_0 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND3_X4 A1 A2 A3 ZN VDD VSS 
M_i_5__m3 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m3 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m3 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m2 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m2 ZN A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m3 VSS A3 net_1__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m3 net_1__m3 A2 net_0__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 net_0__m3 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 ZN A1 net_0__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 net_0__m2 A2 net_1__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m2 net_1__m2 A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 VSS A3 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 net_1__m1 A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 A2 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1__m0_0 A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND3_X2 A1 A2 A3 ZN VDD VSS 
M_i_5__m0_x2__m1 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_x2__m1 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_x2__m1 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_x2__m0 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_x2__m0 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_x2__m0 ZN A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m1 VSS A3 net_1__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_m2__m1 net_1__m0_0__m1 A2 net_0__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m1 net_0__m0_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m0 ZN A1 net_0__m0_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_m2__m0 net_0__m0_0__m0_0 A2 net_1__m0_0__m0_0 VSS NMOS_VTL L=0.050000U 
+ W=0.415000U 
M_i_2__m0_m2__m0 net_1__m0_0__m0_0 A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND2_X2 A1 A2 ZN VDD VSS 
M_i_3__m0_x2__m1 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_x2__m1 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_x2__m0 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_x2__m0 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m0_m2__m1 VSS A2 net_0__m0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m1 net_0__m0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m0 ZN A1 net_0__m0__m0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_m2__m0 net_0__m0__m0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT MUX2_X2 A B S Z VDD VSS 
M_i_11 VDD S x1 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_1_1 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 S Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 Z_neg B net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 net_2 x1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 VDD A net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 VSS S x1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 Z_neg S net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_0 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS x1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 net_1 A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT MUX2_X1 A B S Z VDD VSS 
M_i_1 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD B net_3 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_9 net_3 x1 Z_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_6 net_2 S Z_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_8 VDD A net_2 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_11 VDD S x1 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_0 B VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 Z_neg S net_0 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_5 Z_neg x1 net_1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_4 net_1 A VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_10 VSS S x1 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT LOGIC1_X1 Z VDD VSS 
M_p_tran_2 VDD A Z VDD PMOS_VTL L=0.050000U W=0.135000U 
M_n_tran_1 VSS A A VSS NMOS_VTL L=0.050000U W=0.090000U 
.ENDS

.SUBCKT LOGIC0_X1 Z VDD VSS 
M_transistor_0 VDD A A VDD PMOS_VTL L=0.050000U W=0.090000U 
M_n_tran_1 VSS A Z VSS NMOS_VTL L=0.050000U W=0.090000U 
.ENDS

.SUBCKT INV_X2 A ZN VDD VSS 
M_i_1_0_x2_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x2_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x2_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x2_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT INV_X16 A ZN VDD VSS 
M_i_1_15 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_14 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_13 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_12 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_11 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_10 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_9 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_8 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_7 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_6 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_5 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_4 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_15 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_13 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_12 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_11 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_10 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_9 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_8 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_7 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_6 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_5 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_4 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_3 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT FILLCELL_X8 VDD VSS 
.ENDS

.SUBCKT FILLCELL_X4 VDD VSS 
.ENDS

.SUBCKT FILLCELL_X32 VDD VSS 
.ENDS

.SUBCKT FILLCELL_X2 VDD VSS 
.ENDS

.SUBCKT FILLCELL_X16 VDD VSS 
.ENDS

.SUBCKT FILLCELL_X1 VDD VSS 
.ENDS

.SUBCKT FA_X1 A B CI CO S VDD VSS 
M_instance_315 S net_005 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_instance_275 VDD A net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_280 net_009 B net_010 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_284 net_010 CI net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_290 net_005 net_001 net_011 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_303 net_011 A VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_297 VDD CI net_011 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_309 net_011 B VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_263 VDD B net_008 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_269 net_008 A VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_257 net_001 CI net_008 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_251 net_007 A net_001 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_246 VDD B net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_instance_239 CO net_001 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_instance_233 S net_005 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_instance_194 VSS A net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_199 net_003 B net_004 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_203 net_004 CI net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_209 net_005 net_001 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_221 net_006 A VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_215 VSS CI net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_227 net_006 B VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_182 VSS B net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_188 net_002 A VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_176 net_001 CI net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_170 net_000 A net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_166 VSS B net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_instance_159 CO net_001 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT DLL_X2 D GN Q VDD VSS 
M_i_48 net_000 GN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_92 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_92_11 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_85 VDD net_003 net_005 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_79 VDD net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_73 net_007 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_67 net_003 net_001 net_006 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_62 net_006 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_55 VDD net_000 net_001 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 net_000 GN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_42 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_42_3 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_35 VSS net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_29 VSS net_005 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 VSS net_000 net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DLL_X1 D GN Q VDD VSS 
M_i_48 net_000 GN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_92 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_85 VDD net_003 net_005 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_79 VDD net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_73 net_007 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_67 net_003 net_001 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_62 net_006 D VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_55 VDD net_000 net_001 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 net_000 GN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_42 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_35 VSS net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_29 VSS net_005 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 VSS net_000 net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DLH_X2 D G Q VDD VSS 
M_i_82 VDD net_003 net_005 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_76 VDD net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_72 net_007 net_001 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_66 net_003 net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_61 net_006 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_55 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_89_4 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_89 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_48 VDD G net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_34 VSS net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 VSS net_005 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_000 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_001 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_41_11 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_41 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS G net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DLH_X1 D G Q VDD VSS 
M_i_82 VDD net_003 net_005 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_76 VDD net_005 net_007 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_72 net_007 net_001 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_66 net_003 net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_61 net_006 D VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_55 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_89_4 Q net_003 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_48 VDD G net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_34 VSS net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 VSS net_005 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_000 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_001 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_41_11 Q net_003 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS G net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFF_X2 D CK Q QN VDD VSS 
M_MP13_26 VDD z10 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP13 VDD z10 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP14 QN z9 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP14_5 QN z9 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP10 VDD z9 z10 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP11 z11 z10 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP12 z9 ci z11 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP9 z9 cni z7 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP8 z7 z3 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP1 VDD CK cni VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP5 z4 z3 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP3 z5 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP4 z3 ci z5 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP7 z1 cni z3 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP6 VDD z4 z1 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP2 ci cni VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MN13_38 VSS z10 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN13 VSS z10 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN14 QN z9 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN14_8 QN z9 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN10 VSS z9 z10 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN11 z8 z10 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN12 z9 cni z8 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN9 z9 ci z12 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN8 z12 z3 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN1 VSS CK cni VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN5 z4 z3 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN3 z2 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN4 z2 cni z3 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN7 z3 ci z6 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN6 VSS z4 z6 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN2 ci cni VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFFS_X2 D SN CK Q QN VDD VSS 
M_i_142 VDD net_010 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_189_10 QN net_010 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_189 QN net_010 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_182 VDD net_007 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_182_20 VDD net_007 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_149 net_015 SN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_165 VDD net_007 net_015 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_161 net_015 net_001 net_010 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_176 net_010 net_000 net_016 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_171 net_016 net_003 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_92 VDD CK net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_134 VDD net_003 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_128 net_006 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_122 VDD net_006 net_013 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_118 net_013 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_111 net_003 net_001 net_012 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_106 net_012 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_99 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_46 VSS net_010 net_007 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_86_15 QN net_010 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_86 QN net_010 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_79 VSS net_007 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_79_29 VSS net_007 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_53 net_008 SN VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_59 net_009 net_007 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_63 net_010 net_000 net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_69 net_011 net_001 net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_73 VSS net_003 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS CK net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_006 net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_36 net_005 SN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_30 VSS net_006 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_25 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_19 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_15 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFFS_X1 D SN CK Q QN VDD VSS 
M_i_182 VDD net_007 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_189 QN net_010 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_142 VDD net_010 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_149 net_015 SN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_165 VDD net_007 net_015 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_161 net_015 net_001 net_010 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_176 net_010 net_000 net_016 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_171 net_016 net_003 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_92 VDD CK net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_134 VDD net_003 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_128 net_006 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_122 VDD net_006 net_013 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_118 net_013 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_111 net_003 net_001 net_012 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_106 net_012 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_99 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_79 VSS net_007 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_86 QN net_010 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_46 VSS net_010 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_53 net_008 SN VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_59 net_009 net_007 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_63 net_010 net_000 net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_69 net_011 net_001 net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_73 VSS net_003 net_011 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS CK net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_40 net_006 net_003 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_36 net_005 SN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_30 VSS net_006 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_25 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_19 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_15 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFFR_X2 D RN CK Q QN VDD VSS 
M_i_187_39 Q net_011 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_187 Q net_011 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_180 VDD net_008 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_180_3 VDD net_008 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_172 VDD net_008 net_011 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_165 net_011 RN VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_159 VDD net_011 net_016 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_153 net_016 net_001 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_147 net_008 net_000 net_015 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 net_015 net_003 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_136 VDD net_003 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_125 net_013 RN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_119 VDD net_006 net_013 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_114 net_013 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_108 net_003 net_001 net_012 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_103 net_012 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_96 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_89 VDD CK net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_83_49 Q net_011 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_83 Q net_011 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_76 VSS net_008 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_76_4 VSS net_008 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_70 net_011 net_008 net_010 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_65 net_010 RN VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_59 VSS net_011 net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_55 net_009 net_000 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_49 net_008 net_001 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_45 net_007 net_003 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_38 VSS net_003 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_32 VSS RN net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 net_005 net_006 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS CK net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFFR_X1 D RN CK Q QN VDD VSS 
M_i_187 Q net_011 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_180 VDD net_008 QN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_172 VDD net_008 net_011 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_165 net_011 RN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_159 VDD net_011 net_016 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_153 net_016 net_001 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_147 net_008 net_000 net_015 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_143 net_015 net_003 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_136 VDD net_003 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_125 net_013 RN VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_119 VDD net_006 net_013 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_114 net_013 net_000 net_003 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_108 net_003 net_001 net_012 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_103 net_012 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_96 net_001 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_89 VDD CK net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_83 Q net_011 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_76 VSS net_008 QN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_70 net_011 net_008 net_010 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_65 net_010 RN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_59 VSS net_011 net_009 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_55 net_009 net_000 net_008 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_49 net_008 net_001 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_45 net_007 net_003 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_38 VSS net_003 net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_32 VSS RN net_005 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_28 net_005 net_006 net_004 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_24 net_004 net_001 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_18 net_003 net_000 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_002 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS CK net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT DFFRS_X2 D RN SN CK Q QN VDD VSS 
M_MP91 ckn_i CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP11 VDD D np1 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP12 np1 ck_i z37 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP34 np32 ckn_i z37 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP31 VDD z51 np32 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP33 VDD RN np32 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP101 ck_i ckn_i VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP22 z51 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP21 VDD z37 z51 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP42 VDD z37 np4 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP41 np4 ckn_i z41 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP62 np61 ck_i z41 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP61 VDD z56 np61 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP63 VDD SN np61 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP51 z56 z41 VDD VDD PMOS_VTL L=0.050000U W=0.485000U 
M_MP52 VDD RN z56 VDD PMOS_VTL L=0.050000U W=0.485000U 
M_transistor_3 z99 SN VDD VDD PMOS_VTL L=0.050000U W=0.485000U 
M_transistor_2 VDD z56 z99 VDD PMOS_VTL L=0.050000U W=0.485000U 
M_MP81_1_55 VDD z56 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP81_1 VDD z56 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP81_0 QN z99 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP81_0_51 QN z99 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MN91 ckn_i CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN12 nn1 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN11 z37 ckn_i nn1 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN31 nn31 ck_i z37 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN32 nn32 z51 nn31 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN33 VSS RN nn32 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN101 VSS ckn_i ck_i VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MP91_1 nn2 SN z51 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MP91_0 VSS z37 nn2 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN42 nn4 z37 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN41 z41 ck_i nn4 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN61 nn61 ckn_i z41 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN62 nn62 z56 nn61 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN63 VSS SN nn62 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN52 nn5 z41 z56 VSS NMOS_VTL L=0.050000U W=0.310000U 
M_MN51 VSS RN nn5 VSS NMOS_VTL L=0.050000U W=0.310000U 
M_transistor_1 nn99 SN VSS VSS NMOS_VTL L=0.050000U W=0.310000U 
M_transistor_0 z99 z56 nn99 VSS NMOS_VTL L=0.050000U W=0.310000U 
M_MN91_0_0_58 VSS z56 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN91_0_0 VSS z56 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN81 QN z99 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN81_53 QN z99 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT DFFRS_X1 D RN SN CK Q QN VDD VSS 
M_MP91 ckn_i CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP11 VDD D np1 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP12 np1 ck_i z37 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP34 np32 ckn_i z37 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP31 VDD z51 np32 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP33 VDD RN np32 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP101 ck_i ckn_i VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP22 z51 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP21 VDD z37 z51 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP42 VDD z37 np4 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP41 np4 ckn_i z41 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP62 np61 ck_i z41 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP61 VDD z56 np61 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP63 VDD SN np61 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP52 VDD RN z56 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP51 z56 z41 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_transistor_3 z99 SN VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_transistor_2 VDD z56 z99 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP81_1 VDD z56 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP81_0 QN z99 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MN91 ckn_i CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN12 nn1 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN11 z37 ckn_i nn1 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN31 nn31 ck_i z37 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN32 nn32 z51 nn31 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN33 VSS RN nn32 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN101 VSS ckn_i ck_i VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MP91_1 nn2 SN z51 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MP91_0 VSS z37 nn2 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN42 nn4 z37 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN41 z41 ck_i nn4 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN61 nn61 ckn_i z41 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN62 nn62 z56 nn61 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN63 VSS SN nn62 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN52 nn5 RN z56 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN51 VSS z41 nn5 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_transistor_1 nn99 SN VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_transistor_0 z99 z56 nn99 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN91_0_0 VSS z56 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN81 QN z99 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT CLKGATE_X8 CK E GCK VDD VSS 
M_i_109_4_19_36 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_24_52 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_4_22 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_53 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_4_19 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_24 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_4 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103_74_97 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97_71_87 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97_99 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103_72 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103_74 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97_71 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_90 VDD CK net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_57_165 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_57 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_64 net_008 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_78 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_84 net_004 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_51_7_25_30 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_10_28 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_7_58 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_40 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_7_25 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_10 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_7 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_45_66_78 VSS net_000 net_007d VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40_75_82 net_007d CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40_71 net_007c CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_45_63 VSS net_000 net_007c VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_45_66 VSS net_000 net_007 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40_75 net_007 CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40 net_007b CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_45 VSS net_000 net_007b VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_33 VSS CK net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0_174 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_21 VSS E net_003 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_27 net_004 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATE_X4 CK E GCK VDD VSS 
M_i_109_4_19 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_24 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109_4 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103_74 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97_71 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_90 VDD CK net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_84 net_004 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_64 net_008 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_78 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_57 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_51_7_25 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_10 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51_7 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_45_66 VSS net_000 net_007 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40_75 net_007 CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40 net_007b CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_45 VSS net_000 net_007b VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_33 VSS CK net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 net_004 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_21 VSS E net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT CLKGATE_X2 CK E GCK VDD VSS 
M_i_109_4 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_109 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_103 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_90 VDD CK net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_84 net_004 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_64 net_008 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_78 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_57 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_51_7 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_51 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_45 VSS net_000 net_007 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_40 net_007 CK net_006 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_33 VSS CK net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 net_004 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_21 VSS E net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATE_X1 CK E GCK VDD VSS 
M_i_109 GCK net_006 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_97 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_103 VDD net_000 net_006 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_90 VDD CK net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_84 net_004 net_005 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_78 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_74 net_009 net_004 net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_68 net_002 net_005 net_008 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_64 net_008 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_57 VDD net_002 net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_51 GCK net_006 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_40 net_007 CK net_006 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_45 VSS net_000 net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_33 VSS CK net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 net_004 net_005 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_21 VSS E net_003 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_17 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_11 net_002 net_004 net_001 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_7 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_0 VSS net_002 net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATETST_X8 CK E SE GCK VDD VSS 
M_i_133_10_28_7 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_11_14 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_10_20 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_38 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_10_28 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_11 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_10 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120_72_145 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127_69_164 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127_158 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120_163 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120_72 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127_69 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_114 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_101 net_004 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_101_94 net_004 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_95 VDD net_004 net_011 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_80 net_010 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_107 VDD net_006 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_74 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_69 net_009 SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_63_13_29_4 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_15_27 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_13_55 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_12 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_13_29 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_15 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_13 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_52_76_137 net_008d CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57_77_169 net_007 net_002 net_008d VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57_123 net_007 net_002 net_008c VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_52_150 net_008c CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_52_76 net_008b CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57_77 net_007 net_002 net_008b VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57 net_007 net_002 net_008 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_52 net_008 CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_46 net_006 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_33 net_004 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_33_93 net_004 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_27 VSS net_004 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_39 VSS net_006 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 VSS E net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 net_000 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATETST_X4 CK E SE GCK VDD VSS 
M_i_133_10_28 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_11 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133_10 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120_72 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127_69 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_114 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_101 net_004 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_95 VDD net_004 net_011 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_80 net_010 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_107 VDD net_006 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_74 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_69 net_009 SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_63_13_29 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_15 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63_13 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_52_76 net_008b CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57_77 net_007 net_002 net_008b VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57 net_007 net_002 net_008 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_52 net_008 CK VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_46 net_006 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_33 net_004 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_27 VSS net_004 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_39 VSS net_006 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 VSS E net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 net_000 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATETST_X2 CK E SE GCK VDD VSS 
M_i_114 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_133_10 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_133 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_120 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_101 net_004 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_95 VDD net_004 net_011 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_80 net_010 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_69 net_009 SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_74 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_107 VDD net_006 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_46 net_006 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_63_13 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_63 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_52 net_008 CK net_007 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_57 VSS net_002 net_008 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_33 net_004 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 VSS net_004 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_0 net_000 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 VSS E net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_39 VSS net_006 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKGATETST_X1 CK E SE GCK VDD VSS 
M_i_133 GCK net_007 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_127 VDD net_002 net_007 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_120 net_007 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_114 net_006 CK VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_101 net_004 net_002 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_107 VDD net_006 net_005 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_95 VDD net_004 net_011 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_91 net_011 net_006 net_002 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_i_85 net_002 net_005 net_010 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_80 net_010 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_i_74 VDD E net_009 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_69 net_009 SE net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_63 GCK net_007 VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_57 VSS net_002 net_008 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_52 net_008 CK net_007 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_46 net_006 CK VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_33 net_004 net_002 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_39 VSS net_006 net_005 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_27 VSS net_004 net_003 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_23 net_003 net_005 net_002 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_i_17 net_002 net_006 net_001 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_13 net_001 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_i_7 VSS E net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 net_000 SE VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT CLKBUF_X3 A Z VDD VSS 
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_2_1 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.195000U 
.ENDS

.SUBCKT CLKBUF_X2 A Z VDD VSS 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_2 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.195000U 
.ENDS

.SUBCKT BUF_X8 A Z VDD VSS 
M_i_1_7 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_6 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_5 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_4 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_2 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_0 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_7 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_6 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_5 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_4 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_3 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_2 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT BUF_X4 A Z VDD VSS 
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_0 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT BUF_X2 A Z VDD VSS 
M_i_1_0_x2_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x2_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x2_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x2_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT BUF_X16 A Z VDD VSS 
M_i_1_15 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_14 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_13 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_12 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_11 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_10 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_9 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_8 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_7 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_6 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_5 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_4 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_7 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_6 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_5 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_4 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_2 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_0 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_15 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_13 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_12 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_11 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_10 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_9 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_8 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_7 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_6 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_5 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_4 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_7 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_6 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_5 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_4 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_3 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_2 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI22_X4 A1 A2 B1 B2 ZN VDD VSS 
M_i_5__m3 net_2 A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m3 ZN A1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 net_2 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m2 ZN A2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 net_2 A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 ZN A1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 net_2 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN A2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m3 net_2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m3 VDD B1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m2 net_2 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m2 VDD B2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 net_2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 VDD B1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_2 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD B2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m3 VSS A2 net_0__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 net_0__m3 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 ZN A1 net_0__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 net_0__m2 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 VSS A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m3 VSS B2 net_1__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m3 net_1__m3 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m2 ZN B1 net_1__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m2 net_1__m2 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 VSS B2 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_1__m1 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 ZN B1 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_1__m0_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI22_X2 A1 A2 B1 B2 ZN VDD VSS 
M_i_5__m1 net_2 A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 ZN A1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 net_2 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN A2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 net_2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 VDD B1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_2 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD B2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 VSS A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 VSS B2 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_1__m1 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 ZN B1 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_1__m0_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI222_X4 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_15_3_x4_0 VDD ZN_6 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_1 ZN ZN_6 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_2 VDD ZN_6 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15_3_x4_3 ZN ZN_6 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x2_1 VDD ZN_5 ZN_6 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x2_0 ZN_6 ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11 VDD C2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 net_4 C1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_3 B1 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 net_4 B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_3 A2 ZN_5 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 ZN_5 A1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_14_0_x4_3 VSS ZN_6 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_2 ZN ZN_6 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_1 VSS ZN_6 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_14_0_x4_0 ZN ZN_6 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x2_1 VSS ZN_5 ZN_6 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x2_0 ZN_6 ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS C2 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 net_2 C1 ZN_5 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN_5 B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 A1 ZN_5 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI222_X2 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_7__m0 net_3 A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 ZN A2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_3 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 ZN A1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 net_4 B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 net_3 B1 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 net_4 B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 net_3 B2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11__m1 net_4 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10__m1 VDD C1 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10__m0 net_4 C1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11__m0 VDD C2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m0 net_0__m0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 VSS A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN A1 net_0__m0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS B2 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 net_1__m0_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 ZN B1 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_1__m1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m0 VSS C2 net_2__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 net_2__m0_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 ZN C1 net_2__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m1 net_2__m1 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI221_X4 A B1 B2 C1 C2 ZN VDD VSS 
M_i_13_0_x4_3 VDD ZN_5 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x4_2 ZN ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x4_1 VDD ZN_5 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_13_0_x4_0 ZN ZN_5 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_1_x2_0 VDD ZN_4 ZN_5 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_1_x2_1 ZN_5 ZN_4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 VDD B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_3 A net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 C2 ZN_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 ZN_4 C1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_12_0_x4_3 VSS ZN_5 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_2 ZN ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_1 VSS ZN_5 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_12_0_x4_0 ZN ZN_5 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_0_x2_1 VSS ZN_4 ZN_5 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_0_x2_0 ZN_5 ZN_4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 B1 ZN_4 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN_4 A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 VSS C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 C1 ZN_4 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI221_X2 A B1 B2 C1 C2 ZN VDD VSS 
M_i_6__m1 net_2 C2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN C1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m1 net_2 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 ZN C2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_0 net_2 A net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 net_3 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 VDD B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 net_3 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 VDD B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7_1 net_3 A net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 VSS C2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN C1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 ZN B1 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 net_1__m1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 VSS B2 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_1__m0_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI21_X4 A B1 B2 ZN VDD VSS 
M_i_4__m3 net_1 B2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m3 ZN B1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m2 net_1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m2 ZN B2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 net_1 B2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m1 ZN B1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0 net_1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 ZN B2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_3 net_1 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_2 VDD A net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_1 net_1 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_0 VDD A net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m3 VSS B2 net_0__m3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m3 net_0__m3 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m2 ZN B1 net_0__m2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m2 net_0__m2 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m1 VSS B2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN B1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_3 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_2 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI21_X2 A B1 B2 ZN VDD VSS 
M_i_4__m0_x2__m1 net_1 B2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_x2__m0 ZN B1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_x2__m1 net_1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_x2__m0 ZN B2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_0_x2_1 net_1 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5_0_x2_0 VDD A net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m0_m2__m0 VSS B2 net_0__m0_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m0 net_0__m0_0__m0_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_m2__m1 ZN B1 net_0__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_m2__m1 net_0__m0_0__m1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0_x2_0 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0_x2_1 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI211_X4 A B C1 C2 ZN VDD VSS 
M_i_11_3 VDD ZN_4 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_2 ZN ZN_4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_1 VDD ZN_4 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11_0 ZN ZN_4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9_1 VDD ZN_3 ZN_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9_0 ZN_4 ZN_3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 B net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_1 C2 ZN_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN_3 C1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10_3 VSS ZN_4 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_2 ZN ZN_4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_1 VSS ZN_4 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_10_0 ZN ZN_4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_8_1 VSS ZN_3 ZN_4 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_8_0 ZN_4 ZN_3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A ZN_3 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN_3 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 VSS C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 C1 ZN_3 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI211_X2 A B C1 C2 ZN VDD VSS 
M_i_5__m1 net_1 C2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m1 ZN C1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0 net_1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0 ZN C2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 net_1 B net_2__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 net_2__m1 A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 VDD A net_2__m0_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 net_2__m0_0 B net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m1 VSS C2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m1 net_0__m1 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0 ZN C1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0 net_0__m0_0 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 VSS B ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 ZN B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT ANTENNA_X1 A VDD VSS 
.ENDS

.SUBCKT AND4_X4 A1 A2 A3 A4 ZN VDD VSS 
M_i_1_3 VDD x1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 ZN x1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD x1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN x1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m1 VDD A4 x1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m1 x1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m1 VDD A2 x1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m1 x1 A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0 VDD A1 x1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0 x1 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8__m0 VDD A3 x1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9__m0 x1 A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_3 VSS x1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN x1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS x1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN x1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m1 VSS A4 net_2__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m1 net_2__m1 A3 net_1__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m1 net_1__m1 A2 net_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m1 net_0__m1 A1 x1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0 x1 A1 net_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0 net_0__m0_0 A2 net_1__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0 net_1__m0_0 A3 net_2__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5__m0 net_2__m0_0 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND4_X2 A1 A2 A3 A4 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD A4 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 ZN_neg A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS A4 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 net_2 A3 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND4_X1 A1 A2 A3 A4 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD A4 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_8 ZN_neg A3 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_7 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_6 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS A4 net_2 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_4 net_2 A3 net_1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_3 net_1 A2 net_0 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT AND3_X4 A1 A2 A3 ZN VDD VSS 
M_i_1_0_x4_3 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_2 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0_x2__m1 VDD A3 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0_x2__m1 ZN_neg A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_x2__m1 VDD A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_x2__m0 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6__m0_x2__m0 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7__m0_x2__m0 ZN_neg A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x4_3 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_2 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4__m0_m2__m1 VSS A3 net_1__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_m2__m1 net_1__m0_0__m1 A2 net_0__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_m2__m1 net_0__m0_0__m1 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_m2__m0 ZN_neg A1 net_0__m0_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_m2__m0 net_0__m0_0__m0_0 A2 net_1__m0_0__m0_0 VSS NMOS_VTL L=0.050000U 
+ W=0.415000U 
M_i_4__m0_m2__m0 net_1__m0_0__m0_0 A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND3_X2 A1 A2 A3 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A3 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 ZN_neg A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 VDD A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS A3 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND2_X4 A1 A2 ZN VDD VSS 
M_i_1_0_x4_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_2 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_0 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_3 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_x2__m0 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_x2__m1 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4__m0_x2__m0 VDD A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5__m0_x2__m1 ZN_neg A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x4_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_2 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_3 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_m2__m1 VSS A2 net_0__m0_0__m1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_m2__m1 net_0__m0_0__m1 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2__m0_m2__m0 ZN_neg A1 net_0__m0_0__m0_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3__m0_m2__m0 net_0__m0_0__m0_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND2_X2 A1 A2 ZN VDD VSS 
M_i_1_1 VDD ZN_neg ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_1 VSS ZN_neg ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT BUF_X32 A Z VDD VSS 
M_i_1_31 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_30 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_29 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_28 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_27 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_26 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_25 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_24 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_23 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_22 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_21 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_20 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_19 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_18 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_17 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_16 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_15 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_14 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_13 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_12 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_11 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_10 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_9 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_8 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_7 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_6 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_5 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_4 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_3 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD Z_neg Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_15 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_14 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_13 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_12 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_11 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_10 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_9 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_8 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_7 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_6 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_5 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_4 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_2 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_0 Z_neg A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_31 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_30 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_29 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_28 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_27 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_26 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_25 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_24 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_23 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_22 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_21 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_20 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_19 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_18 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_17 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_16 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_13 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_12 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_11 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_10 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_9 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_8 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_7 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_6 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_5 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_4 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_3 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS Z_neg Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_15 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_14 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_13 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_12 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_11 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_10 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_9 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_8 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_7 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_6 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_5 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_4 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_3 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_2 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_1 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2_0 Z_neg A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT INV_X8 A ZN VDD VSS 
M_i_1_0_x8_7 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_6 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_5 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_4 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x8_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x8_7 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_6 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_5 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_4 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_3 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_2 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x8_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT INV_X4 A ZN VDD VSS 
M_i_1_0_x4_3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0_x4_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_0_x4_3 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_2 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0_x4_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT CLKBUF_X1 A Z VDD VSS 
M_i_1 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.195000U 
M_i_2 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.095000U 
.ENDS

.SUBCKT INV_X32 A ZN VDD VSS 
M_i_1_31 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_30 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_29 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_28 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_27 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_26 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_25 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_24 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_23 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_22 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_21 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_20 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_19 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_18 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_17 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_16 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_15 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_14 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_13 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_12 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_11 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_10 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_9 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_8 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_7 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_6 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_5 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_4 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_3 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_2 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_1 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1_0 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_31 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_30 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_29 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_28 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_27 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_26 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_25 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_24 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_23 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_22 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_21 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_20 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_19 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_18 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_17 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_16 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_15 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_14 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_13 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_12 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_11 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_10 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_9 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_8 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_7 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_6 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_5 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_4 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_3 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI221_X1 A B1 B2 C1 C2 ZN VDD VSS 
M_i_5 net_2 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 ZN C2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 A net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_3 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD B2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 ZN B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 net_1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT DFF_X1 D CK Q QN VDD VSS 
M_MP13 VDD z10 Q VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP14 QN z9 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_MP10 VDD z9 z10 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP11 z11 z10 VDD VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP12 z9 ci z11 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP9 z9 cni z7 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP8 z7 z3 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP1 VDD CK cni VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP5 z4 z3 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MP3 z5 D VDD VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP4 z3 ci z5 VDD PMOS_VTL L=0.050000U W=0.420000U 
M_MP7 z1 cni z3 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP6 VDD z4 z1 VDD PMOS_VTL L=0.050000U W=0.090000U 
M_MP2 ci cni VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_MN13 VSS z10 Q VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN14 QN z9 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_MN10 VSS z9 z10 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN11 z8 z10 VSS VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN12 z9 cni z8 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN9 z9 ci z12 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN8 z12 z3 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN1 VSS CK cni VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN5 z4 z3 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_MN3 z2 D VSS VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN4 z2 cni z3 VSS NMOS_VTL L=0.050000U W=0.275000U 
M_MN7 z3 ci z6 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN6 VSS z4 z6 VSS NMOS_VTL L=0.050000U W=0.090000U 
M_MN2 ci cni VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT OR3_X1 A1 A2 A3 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A3 net_1 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_6 net_1 A2 net_0 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_5 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS A3 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_3 ZN_neg A2 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 VSS A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT OR4_X1 A1 A2 A3 A4 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 VDD A4 net_2 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_8 net_2 A3 net_1 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_7 net_1 A2 net_0 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_6 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS A4 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_4 ZN_neg A3 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT AOI211_X1 A B C1 C2 ZN VDD VSS 
M_i_7 VDD A net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 B net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_1 C1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 ZN C2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS B ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN C1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI222_X1 A1 A2 B1 B2 C1 C2 ZN VDD VSS 
M_i_6 net_3 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 ZN A2 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_9 net_3 B2 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_8 net_4 B1 net_3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 VDD C1 net_4 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_11 net_4 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS B2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 ZN C1 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 net_2 C2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI22_X1 A1 A2 B1 B2 ZN VDD VSS 
M_i_5 VDD A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 ZN B1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 net_2 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1 net_0 A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_0 B1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT XNOR2_X1 A B ZN VDD VSS 
M_i_53 VDD B net_003 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_48 net_003 A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_42 ZN net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_36 VDD B net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_29 net_000 A VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_23 net_002 B ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_17 ZN A net_002 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_11 net_002 net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_5 VSS B net_001 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 net_001 A net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT AOI21_X1 A B1 B2 ZN VDD VSS 
M_i_5 VDD A net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 net_1 B1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN B2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2 VSS A ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 ZN B1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI211_X1 A B C1 C2 ZN VDD VSS 
M_i_7 ZN B VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN C1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_2 C2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 VSS B net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 C1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN C2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AOI22_X1 A1 A2 B1 B2 ZN VDD VSS 
M_i_5 net_2 A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 ZN A1 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 net_2 B1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD B2 net_2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN B1 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_1 B2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND2_X1 A1 A2 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 VDD A2 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_4 ZN_neg A1 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT NAND2_X1 A1 A2 ZN VDD VSS 
M_i_2 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT AND3_X1 A1 A2 A3 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 VDD A3 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_6 ZN_neg A2 VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_5 VDD A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_4 VSS A3 net_1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_3 net_1 A2 net_0 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 net_0 A1 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT NAND4_X1 A1 A2 A3 A4 ZN VDD VSS 
M_i_4 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_6 VDD A3 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_7 ZN A4 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 A3 net_2 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 net_2 A4 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR2_X1 A1 A2 ZN VDD VSS 
M_i_2 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 net_0 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OAI21_X1 A B1 B2 ZN VDD VSS 
M_i_5 VDD A ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 ZN B1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_1 B2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2 VSS A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 net_0 B1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 ZN B2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND3_X1 A1 A2 A3 ZN VDD VSS 
M_i_3 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 ZN A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 A2 net_1 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 net_1 A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NOR3_X1 A1 A2 A3 ZN VDD VSS 
M_i_3 ZN A1 net_0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 net_0 A2 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 net_1 A3 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 ZN A3 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT OR2_X1 A1 A2 ZN VDD VSS 
M_i_1 ZN ZN_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_5 VDD A2 net_0 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_4 net_0 A1 ZN_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 ZN ZN_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_3 VSS A2 ZN_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 ZN_neg A1 VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT NOR2_X4 A1 A2 ZN VDD VSS 
M_i_3__m0_m2__m1 VDD A2 net_0__m0__m1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m1 net_0__m0__m1 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m0 ZN A1 net_0__m0__m0 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_m2__m0 net_0__m0__m0 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_m2__m1_58 VDD A2 net_0__m0__m2 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m1_45 net_0__m0__m2 A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2__m0_m2__m0_52 ZN A1 net_0__m0__m3 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3__m0_m2__m0_38 net_0__m0__m3 A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_1__m0_x2__m1 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m1 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m0 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_x2__m0 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_x2__m1_23 VSS A2 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m1_57 ZN A1 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0__m0_x2__m0_35 VSS A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1__m0_x2__m0_16 ZN A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT NAND2_X4 A1 A2 ZN VDD VSS 
M_i_2_3 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_2 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_1 VDD A1 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_2_0 ZN A1 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_3 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_2 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_1 VDD A2 ZN VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3_0 ZN A2 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0_3 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_2 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_1 net_0 A1 ZN VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0_0 ZN A1 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_3 net_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_2 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_1 net_0 A2 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1_0 VSS A2 net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT BUF_X1 A Z VDD VSS 
M_i_1 Z Z_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 VDD A Z_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_0 Z Z_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_2 VSS A Z_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT HA_X1 A B CO S VDD VSS 
M_i_11 CO CO_neg VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_15 VDD B CO_neg VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_14 CO_neg A VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_8 x1 A net_2 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_9 net_2 B VDD VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_5 VDD x1 net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_3 net_1 A S VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_4 S B net_1 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_10 CO CO_neg VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_13 VSS B net_3 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_12 net_3 A CO_neg VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_6 VSS A x1 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_7 x1 B VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_2 VSS x1 S VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_0 S A net_0 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_1 net_0 B VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT INV_X1 A ZN VDD VSS 
M_i_1 ZN A VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_0 ZN A VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
.ENDS

.SUBCKT XOR2_X1 A B Z VDD VSS 
M_i_53 net_003 B Z VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_47 Z A net_003 VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_41 net_003 net_000 VDD VDD PMOS_VTL L=0.050000U W=0.630000U 
M_i_35 VDD B net_002 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_30 net_002 A net_000 VDD PMOS_VTL L=0.050000U W=0.315000U 
M_i_24 VSS B net_001 VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_19 net_001 A Z VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_13 Z net_000 VSS VSS NMOS_VTL L=0.050000U W=0.415000U 
M_i_7 VSS B net_000 VSS NMOS_VTL L=0.050000U W=0.210000U 
M_i_0 net_000 A VSS VSS NMOS_VTL L=0.050000U W=0.210000U 
.ENDS

.SUBCKT cruisecontrol_DW01_inc_0 SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] 
+ SUM[0] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] VDD VSS 
XU1_1_6 A[6] carry[6] carry[7] SUM[6] VDD VSS HA_X1 
XU1_1_5 A[5] carry[5] carry[6] SUM[5] VDD VSS HA_X1 
XU1_1_4 A[4] carry[4] carry[5] SUM[4] VDD VSS HA_X1 
XU1_1_3 A[3] carry[3] carry[4] SUM[3] VDD VSS HA_X1 
XU1_1_2 A[2] carry[2] carry[3] SUM[2] VDD VSS HA_X1 
XU1_1_1 A[1] A[0] carry[2] SUM[1] VDD VSS HA_X1 
XU1 A[0] SUM[0] VDD VSS INV_X1 
XU2 carry[7] A[7] SUM[7] VDD VSS XOR2_X1 
.ENDS

.SUBCKT cruisecontrol_DW01_inc_1 SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] 
+ SUM[0] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] VDD VSS 
XU1_1_6 A[6] carry[6] carry[7] SUM[6] VDD VSS HA_X1 
XU1_1_5 A[5] carry[5] carry[6] SUM[5] VDD VSS HA_X1 
XU1_1_4 A[4] carry[4] carry[5] SUM[4] VDD VSS HA_X1 
XU1_1_3 A[3] carry[3] carry[4] SUM[3] VDD VSS HA_X1 
XU1_1_2 A[2] carry[2] carry[3] SUM[2] VDD VSS HA_X1 
XU1_1_1 A[1] A[0] carry[2] SUM[1] VDD VSS HA_X1 
XU1 A[0] SUM[0] VDD VSS INV_X1 
XU2 carry[7] A[7] SUM[7] VDD VSS XOR2_X1 
.ENDS

.SUBCKT cruisecontrol speed[7] speed[6] speed[5] speed[4] speed[3] speed[2] speed[1] 
+ speed[0] cruisespeed[7] cruisespeed[6] cruisespeed[5] cruisespeed[4] cruisespeed[3] 
+ cruisespeed[2] cruisespeed[1] cruisespeed[0] reset clk cruisectrl brake resume 
+ cancel coast accel set throttle 
XU71 n300 n295 VDD VSS INV_X1 
XU70 n293 n294 VDD VSS INV_X32 
XU69 n136 n293 VDD VSS INV_X1 
XU68 n290 n292 VDD VSS INV_X32 
XU67 n294 n291 VDD VSS INV_X1 
XU66 n291 n290 VDD VSS CLKBUF_X1 
XU65 n287 n289 VDD VSS INV_X32 
XU64 n1350 n288 VDD VSS INV_X1 
XU63 n286 n287 VDD VSS INV_X1 
XU62 n288 n286 VDD VSS INV_X32 
XU61 n289 n285 VDD VSS BUF_X1 
XU60 n283 n284 VDD VSS INV_X32 
XU59 n137 n283 VDD VSS INV_X1 
XU58 n280 n282 VDD VSS INV_X32 
XU57 n284 n281 VDD VSS INV_X1 
XU56 n281 n280 VDD VSS CLKBUF_X1 
XU55 n278 n279 VDD VSS INV_X32 
XU54 n1340 n278 VDD VSS INV_X1 
XU53 n275 n277 VDD VSS INV_X32 
XU52 n279 n276 VDD VSS INV_X1 
XU51 n276 n275 VDD VSS CLKBUF_X1 
XU50 n270 n274 VDD VSS INV_X32 
XU49 n272 n273 VDD VSS INV_X1 
XU48 n271 n272 VDD VSS INV_X32 
XU47 n1470 n271 VDD VSS INV_X1 
XU46 n273 n270 VDD VSS CLKBUF_X1 
XU45 n265 n269 VDD VSS INV_X32 
XU44 n267 n268 VDD VSS INV_X1 
XU43 n266 n267 VDD VSS INV_X32 
XU42 n1330 n266 VDD VSS INV_X1 
XU41 n268 n265 VDD VSS CLKBUF_X1 
XU40 n260 n264 VDD VSS INV_X32 
XU39 n262 n263 VDD VSS INV_X1 
XU38 n261 n262 VDD VSS INV_X32 
XU37 n1320 n261 VDD VSS INV_X1 
XU36 n263 n260 VDD VSS CLKBUF_X1 
XU35 n255 n259 VDD VSS INV_X32 
XU34 n257 n258 VDD VSS INV_X1 
XU33 n256 n257 VDD VSS INV_X32 
XU32 n1310 n256 VDD VSS INV_X1 
XU31 n258 n255 VDD VSS CLKBUF_X1 
XU30 n253 n254 VDD VSS INV_X32 
XU29 n1300 n253 VDD VSS INV_X1 
XU28 n250 n252 VDD VSS INV_X32 
XU27 n254 n251 VDD VSS INV_X1 
XU26 n251 n250 VDD VSS CLKBUF_X1 
XU25 n129 n249 VDD VSS BUF_X32 
XU24 n246 n248 VDD VSS INV_X32 
XU23 n249 n247 VDD VSS INV_X1 
XU22 n247 n246 VDD VSS CLKBUF_X1 
XU21 n241 n245 VDD VSS INV_X32 
XU20 n243 n244 VDD VSS INV_X1 
XU19 n242 n243 VDD VSS INV_X32 
XU18 n1280 n242 VDD VSS INV_X1 
XU17 n244 n241 VDD VSS CLKBUF_X1 
XU16 n190 n240 VDD VSS INV_X32 
XU15 n1460 n239 VDD VSS INV_X1 
XU14 n235 n238 VDD VSS INV_X1 
XU13 n239 n235 VDD VSS INV_X32 
XU12 n238 n190 VDD VSS CLKBUF_X1 
XU11 n330 n189 VDD VSS BUF_X1 
XU10 n325 n170 VDD VSS BUF_X1 
XU9 n319 n169 VDD VSS BUF_X1 
XU8 n316 n168 VDD VSS BUF_X1 
XU7 n303 n167 VDD VSS BUF_X1 
XU6 n292 n166 VDD VSS BUF_X1 
XU5 n282 n165 VDD VSS BUF_X1 
XU4 n153 n164 VDD VSS INV_X8 
XU3 n277 n153 VDD VSS INV_X1 
XU2 n296 n152 VDD VSS BUF_X1 
XU1 n81 n1 VDD VSS INV_X1 
XINV_X1_G1B2I1 clk clk_G1B7I1 VDD VSS INV_X4 
XINV_X1_G1B1I2 clk_G1B7I1 clk_G1B8I2 VDD VSS INV_X4 
XINV_X1_G1B1I3 clk_G1B7I1 clk_G1B8I3 VDD VSS INV_X4 
XINV_X1_G1B1I1 clk_G1B7I1 clk_G1B8I1 VDD VSS INV_X4 
XU113 n336 n337 VDD VSS INV_X32 
XU112 n143 n336 VDD VSS INV_X1 
XU111 n333 n335 VDD VSS INV_X32 
XU110 n337 n334 VDD VSS INV_X1 
XU109 n334 n333 VDD VSS CLKBUF_X1 
XU108 n331 n332 VDD VSS INV_X32 
XU107 n142 n331 VDD VSS INV_X1 
XU106 n328 n330 VDD VSS INV_X32 
XU105 n332 n329 VDD VSS INV_X1 
XU104 n329 n328 VDD VSS CLKBUF_X1 
XU103 n326 n327 VDD VSS INV_X1 
XU102 n154 n326 VDD VSS INV_X32 
XU101 n324 n325 VDD VSS INV_X32 
XU100 n323 n324 VDD VSS INV_X1 
XU99 n322 n323 VDD VSS INV_X32 
XU98 n141 n322 VDD VSS INV_X1 
XU97 n320 n321 VDD VSS INV_X32 
XU96 n140 n320 VDD VSS INV_X1 
XU95 n317 n319 VDD VSS INV_X32 
XU94 n321 n318 VDD VSS INV_X1 
XU93 n318 n317 VDD VSS CLKBUF_X1 
XU92 n314 n316 VDD VSS INV_X32 
XU91 n139 n315 VDD VSS INV_X1 
XU90 n313 n314 VDD VSS INV_X1 
XU89 n312 n313 VDD VSS INV_X32 
XU88 n315 n312 VDD VSS CLKBUF_X1 
XU87 n310 n311 VDD VSS INV_X1 
XU86 n215 n310 VDD VSS INV_X32 
XU85 n308 n309 VDD VSS INV_X32 
XU84 n138 n308 VDD VSS INV_X1 
XU83 n306 n307 VDD VSS INV_X32 
XU82 n309 n306 VDD VSS INV_X1 
XU81 n304 n305 VDD VSS INV_X32 
XU80 n144 n304 VDD VSS INV_X1 
XU79 n301 n303 VDD VSS INV_X32 
XU78 n305 n302 VDD VSS INV_X1 
XU77 n302 n301 VDD VSS CLKBUF_X1 
XU76 n299 n300 VDD VSS INV_X32 
XU75 n145 n299 VDD VSS INV_X1 
XU74 n297 n298 VDD VSS INV_X1 
XU73 n216 n297 VDD VSS INV_X32 
XU72 n295 n296 VDD VSS INV_X32 
XU158 n1520 n160 VDD VSS INV_X1 
XU157 n720 n1 n113 VDD VSS NAND2_X1 
XU156 n195 n212 VDD VSS INV_X1 
XU154 n110 n230 VDD VSS INV_X1 
XU153 n81 n79 n80 n78 VDD VSS OAI21_X1 
XU152 n78 n228 VDD VSS INV_X1 
XU151 n79 n81 N189 n101 VDD VSS AND3_X1 
XU150 n231 n229 n114 n79 VDD VSS AND3_X1 
XU149 n740 n223 n68 VDD VSS NAND2_X1 
XU148 n229 n108 n710 VDD VSS NOR2_X1 
XU147 n64 n84 n116 VDD VSS NOR2_X1 
XU146 n106 n229 n117 VDD VSS OR2_X1 
XU145 n116 n117 n700 n223 n86 VDD VSS NAND4_X1 
XU144 n720 n233 n700 n229 n107 VDD VSS OAI22_X1 
XU143 n710 n108 n105 VDD VSS NOR2_X1 
XU142 n107 n226 VDD VSS INV_X1 
XU141 n106 n226 n105 n236 n760 VDD VSS OAI211_X1 
XU140 n1 n127 n84 VDD VSS NOR2_X1 
XU139 n102 n125 n50 VDD VSS AND2_X1 
XU138 n109 n125 n51 VDD VSS AND2_X1 
XU137 n66 n115 n1 n126 VDD VSS OAI21_X1 
XU136 n126 n224 VDD VSS INV_X1 
XU135 n109 n230 n79 n188 n104 VDD VSS AOI211_X1 
XU134 n760 n225 VDD VSS INV_X1 
XU133 n225 n104 n1 n89 VDD VSS OAI21_X1 
XU132 n115 n110 n80 VDD VSS NAND2_X1 
XU131 n109 n102 n115 VDD VSS NOR2_X1 
XU130 n222 n223 n88 VDD VSS NAND2_X1 
XU129 n101 n81 n80 N190 n113 n112 VDD VSS AOI221_X1 
XU128 n112 n227 VDD VSS INV_X1 
XU127 n86 n227 n233 n83 n111 VDD VSS AOI211_X1 
XU126 n111 n222 VDD VSS INV_X1 
XU125 n1 n234 resume n720 n90 VDD VSS OAI22_X1 
XU124 n39 state[2] n38 n81 VDD VSS NOR3_X1 
Xspeed_reg_1_ n335 clk_G1B8I3 speed[1] n210 VDD VSS DFF_X1 
Xspeed_reg_2_ n189 clk_G1B8I3 speed[2] n211 VDD VSS DFF_X1 
Xspeed_reg_3_ n170 clk_G1B8I3 speed[3] n154 VDD VSS DFF_X1 
Xspeed_reg_4_ n169 clk_G1B8I2 speed[4] n213 VDD VSS DFF_X1 
Xspeed_reg_5_ n168 clk_G1B8I2 speed[5] n155 VDD VSS DFF_X1 
Xspeed_reg_6_ n307 clk_G1B8I2 speed[6] n215 VDD VSS DFF_X1 
Xspeed_reg_0_ n167 clk_G1B8I3 speed[0] N70 VDD VSS DFF_X1 
Xspeed_reg_7_ n152 clk_G1B8I1 speed[7] n216 VDD VSS DFF_X1 
Xstate_reg_0_ n166 clk_G1B8I2 state[0] n39 VDD VSS DFF_X1 
Xstate_reg_1_ n338 clk_G1B8I2 state[1] n38 VDD VSS DFF_X1 
Xstate_reg_2_ n165 clk_G1B8I2 state[2] n33 VDD VSS DFF_X1 
Xcruisectrl_reg n164 clk_G1B8I2 cruisectrl n18 VDD VSS DFF_X1 
Xcruisespeed_reg_0_ n274 clk_G1B8I1 cruisespeed[0] n218 VDD VSS DFF_X1 
Xcruisespeed_reg_1_ n269 clk_G1B8I1 cruisespeed[1] n1680 VDD VSS DFF_X1 
Xcruisespeed_reg_2_ n264 clk_G1B8I3 cruisespeed[2] n1690 VDD VSS DFF_X1 
Xcruisespeed_reg_3_ n259 clk_G1B8I3 cruisespeed[3] n209 VDD VSS DFF_X1 
Xcruisespeed_reg_4_ n252 clk_G1B8I3 cruisespeed[4] n1670 VDD VSS DFF_X1 
Xcruisespeed_reg_5_ n248 clk_G1B8I1 cruisespeed[5] n208 VDD VSS DFF_X1 
Xcruisespeed_reg_6_ n245 clk_G1B8I1 cruisespeed[6] n217 VDD VSS DFF_X1 
Xcruisespeed_reg_7_ n240 clk_G1B8I1 cruisespeed[7] NETTRAN_DUMMY_1 VDD VSS DFF_X1 
XU251 n188 N189 VDD VSS INV_X1 
XU250 coast n231 VDD VSS INV_X1 
XU249 throttle n700 n710 n236 n69 VDD VSS OAI22_X1 
XU248 n69 n228 resume n65 n67 VDD VSS AOI211_X1 
XU247 n67 n68 n1350 VDD VSS NOR2_X1 
XU246 brake n234 VDD VSS INV_X1 
XU245 n65 n237 VDD VSS INV_X1 
XU244 n66 n237 n233 n62 VDD VSS OAI21_X1 
XU243 n62 n223 n64 n65 n63 VDD VSS OAI211_X1 
XU242 n63 n62 n18 n1340 VDD VSS OAI21_X1 
XU241 accel n127 n109 VDD VSS AND2_X1 
XU240 n81 n234 cancel n103 VDD VSS NAND3_X1 
XU239 n730 n103 n770 VDD VSS NAND2_X1 
XU238 throttle n229 VDD VSS INV_X1 
XU237 cruisespeed[4] n224 n54 VDD VSS NAND2_X1 
XU236 N167 n50 N150 n51 n55 VDD VSS AOI22_X1 
XU235 n54 n55 n47 n213 n1300 VDD VSS OAI211_X1 
XU234 cruisespeed[0] n224 n123 VDD VSS NAND2_X1 
XU233 n218 n50 N146 n51 n124 VDD VSS AOI22_X1 
XU232 n123 n124 n47 N70 n1470 VDD VSS OAI211_X1 
XU231 cruisespeed[1] n224 n60 VDD VSS NAND2_X1 
XU230 N164 n50 N147 n51 n61 VDD VSS AOI22_X1 
XU229 n60 n61 n47 n210 n1330 VDD VSS OAI211_X1 
XU228 cruisespeed[5] n224 n52 VDD VSS NAND2_X1 
XU227 N168 n50 N151 n51 n53 VDD VSS AOI22_X1 
XU226 n52 n53 n47 n155 n129 VDD VSS OAI211_X1 
XU225 cruisespeed[6] n224 n48 VDD VSS NAND2_X1 
XU224 N169 n50 N152 n51 n49 VDD VSS AOI22_X1 
XU223 n48 n49 n47 n311 n1280 VDD VSS OAI211_X1 
XU222 cruisespeed[2] n224 n580 VDD VSS NAND2_X1 
XU221 N165 n50 N148 n51 n59 VDD VSS AOI22_X1 
XU220 n580 n59 n47 n211 n1320 VDD VSS OAI211_X1 
XU219 cruisespeed[3] n224 n56 VDD VSS NAND2_X1 
XU218 N166 n50 N149 n51 n57 VDD VSS AOI22_X1 
XU217 n56 n57 n47 n327 n1310 VDD VSS OAI211_X1 
XU216 cruisespeed[7] n224 n121 VDD VSS NAND2_X1 
XU215 N170 n50 N153 n51 n122 VDD VSS AOI22_X1 
XU214 n121 n122 n47 n298 n1460 VDD VSS OAI211_X1 
XU213 n1 reset n125 VDD VSS NOR2_X1 
XU212 n84 n83 n233 n82 VDD VSS AOI21_X1 
XU211 n33 n740 n82 n68 n137 VDD VSS OAI22_X1 
XU210 set N58 throttle n108 VDD VSS AND3_X1 
XU209 n760 n228 n770 n750 VDD VSS NOR3_X1 
XU208 n39 n740 n750 n68 n136 VDD VSS OAI22_X1 
XU207 n114 n231 throttle n110 VDD VSS NAND3_X1 
XU206 reset n223 VDD VSS INV_X1 
XU205 n224 reset n116 n47 VDD VSS OR3_X1 
XU204 resume n233 VDD VSS INV_X1 
XU203 n102 n81 n99 VDD VSS AND2_X1 
XU202 throttle n700 n236 n100 VDD VSS AOI21_X1 
XU201 n770 n99 n100 n101 n91 VDD VSS OR4_X1 
XU200 n86 n83 n85 VDD VSS NOR2_X1 
XU199 n38 n85 n233 n730 n740 VDD VSS OAI211_X1 
XU198 n84 reset n64 n108 n66 VDD VSS AOI211_X1 
XU197 coast n114 n102 VDD VSS AND2_X1 
XU196 speed[7] r116_carry[7] N135 VDD VSS XNOR2_X1 
XU195 n2 n89 N135 n90 N77 n91 n98 VDD VSS AOI222_X1 
XU194 n222 n298 n98 n88 n145 VDD VSS OAI22_X1 
XU193 n9 n89 speed[0] n90 N70 n91 n97 VDD VSS AOI222_X1 
XU192 n222 N70 n97 n88 n144 VDD VSS OAI22_X1 
XU191 speed[6] r116_carry[6] N134 VDD VSS XNOR2_X1 
XU190 n3 n89 N134 n90 N76 n91 n87 VDD VSS AOI222_X1 
XU189 n311 n222 n87 n88 n138 VDD VSS OAI22_X1 
XU188 speed[5] r116_carry[5] N133 VDD VSS XNOR2_X1 
XU187 n4 n89 N133 n90 N75 n91 n92 VDD VSS AOI222_X1 
XU186 n155 n222 n92 n88 n139 VDD VSS OAI22_X1 
XU185 speed[4] r116_carry[4] N132 VDD VSS XNOR2_X1 
XU184 n5 n89 N132 n90 N74 n91 n93 VDD VSS AOI222_X1 
XU183 n213 n222 n93 n88 n140 VDD VSS OAI22_X1 
XU182 speed[3] r116_carry[3] N131 VDD VSS XNOR2_X1 
XU181 n6 n89 N131 n90 N73 n91 n94 VDD VSS AOI222_X1 
XU180 n327 n222 n94 n88 n141 VDD VSS OAI22_X1 
XU179 speed[2] speed[1] N130 VDD VSS XNOR2_X1 
XU178 n7 n89 N130 n90 N72 n91 n95 VDD VSS AOI222_X1 
XU177 n211 n222 n95 n88 n142 VDD VSS OAI22_X1 
XU176 n8 n89 n210 n90 N71 n91 n96 VDD VSS AOI222_X1 
XU175 n210 n222 n96 n88 n143 VDD VSS OAI22_X1 
XU174 n127 n232 VDD VSS INV_X1 
XU173 n232 accel n114 VDD VSS NOR2_X1 
XU172 cancel brake n127 VDD VSS NOR2_X1 
XU171 n720 n730 n65 VDD VSS NAND2_X1 
XU170 n64 n236 VDD VSS INV_X1 
XU169 n197 n219 VDD VSS INV_X1 
XU168 n200 n214 VDD VSS INV_X1 
XU167 n163 n172 VDD VSS INV_X1 
XU166 n162 n171 VDD VSS INV_X1 
XU165 n1640 n173 VDD VSS INV_X1 
XU164 n1490 n157 VDD VSS INV_X1 
XU163 n1500 n158 VDD VSS INV_X1 
XU162 n1510 n159 VDD VSS INV_X1 
XU161 n161 n1700 VDD VSS INV_X1 
XU160 n1480 n156 VDD VSS INV_X1 
XU159 n1650 n174 VDD VSS INV_X1 
XU328 n205 n207 n206 N190 VDD VSS OAI21_X1 
XU327 cruisespeed[6] n311 n204 n203 n206 VDD VSS AOI22_X1 
XU326 n201 n202 n214 n204 VDD VSS AOI21_X1 
XU325 n198 n219 n199 n202 VDD VSS AOI21_X1 
XU324 n194 n196 n195 n197 VDD VSS OAI21_X1 
XU323 n191 n193 n192 n196 VDD VSS OAI21_X1 
XU322 n1900 cruisespeed[1] n210 n1890 n193 VDD VSS OAI22_X1 
XU321 n1890 n210 n1900 VDD VSS AND2_X1 
XU320 n218 speed[0] n1890 VDD VSS NOR2_X1 
XU319 n207 n205 n221 n188 VDD VSS AOI21_X1 
XU318 n298 cruisespeed[7] n207 VDD VSS NOR2_X1 
XU317 speed[6] n217 n186 n203 n187 VDD VSS AOI22_X1 
XU316 speed[6] cruisespeed[6] n203 VDD VSS XNOR2_X1 
XU315 n200 n185 n184 n186 VDD VSS AOI21_X1 
XU314 n208 speed[5] n200 VDD VSS NOR2_X1 
XU313 n183 n212 n199 n184 VDD VSS NAND3_X1 
XU312 n182 n198 n199 VDD VSS NOR2_X1 
XU311 cruisespeed[4] n213 n198 VDD VSS AND2_X1 
XU310 n209 speed[3] n195 VDD VSS NOR2_X1 
XU309 n194 n181 n192 n220 n183 VDD VSS OAI211_X1 
XU308 speed[3] n209 n194 VDD VSS NAND2_X1 
XU307 n210 n179 n178 cruisespeed[1] n180 VDD VSS AOI22_X1 
XU306 n210 n179 n178 VDD VSS OR2_X1 
XU305 speed[0] n218 n179 VDD VSS NAND2_X1 
XU304 n181 n191 n192 VDD VSS NAND2_X1 
XU303 cruisespeed[2] n211 n191 VDD VSS NAND2_X1 
XU302 n211 cruisespeed[2] n181 VDD VSS OR2_X1 
XU301 n182 n201 n185 VDD VSS NOR2_X1 
XU300 speed[5] n208 n201 VDD VSS AND2_X1 
XU299 n213 cruisespeed[4] n182 VDD VSS NOR2_X1 
XU298 cruisespeed[7] n298 n205 VDD VSS NAND2_X1 
XU297 n177 n176 N58 VDD VSS NAND2_X1 
XU296 speed[5] n175 speed[4] n176 VDD VSS OAI21_X1 
XU295 speed[3] speed[2] speed[1] n175 VDD VSS AND3_X1 
XU294 speed[7] speed[6] n177 VDD VSS NOR2_X1 
XU293 cruisespeed[7] n1660 N170 VDD VSS XOR2_X1 
XU292 cruisespeed[6] n174 n1660 VDD VSS NOR2_X1 
XU291 cruisespeed[6] n1650 N169 VDD VSS XOR2_X1 
XU290 n174 n1640 n208 N168 VDD VSS OAI21_X1 
XU289 n173 cruisespeed[5] n1650 VDD VSS NOR2_X1 
XU288 n173 n163 n1670 N167 VDD VSS OAI21_X1 
XU287 n172 cruisespeed[4] n1640 VDD VSS NOR2_X1 
XU286 n172 n162 n209 N166 VDD VSS OAI21_X1 
XU285 n171 cruisespeed[3] n163 VDD VSS NOR2_X1 
XU284 n171 n161 n1690 N165 VDD VSS OAI21_X1 
XU283 n1700 cruisespeed[2] n162 VDD VSS NOR2_X1 
XU282 n1700 n218 n1680 N164 VDD VSS OAI21_X1 
XU281 cruisespeed[1] cruisespeed[0] n161 VDD VSS NOR2_X1 
XU280 speed[7] n1530 N77 VDD VSS XOR2_X1 
XU279 speed[6] n160 n1530 VDD VSS NOR2_X1 
XU278 speed[6] n1520 N76 VDD VSS XOR2_X1 
XU277 n160 n1510 n155 N75 VDD VSS OAI21_X1 
XU276 n159 speed[5] n1520 VDD VSS NOR2_X1 
XU275 n159 n1500 n213 N74 VDD VSS OAI21_X1 
XU274 n158 speed[4] n1510 VDD VSS NOR2_X1 
XU273 n158 n1490 n327 N73 VDD VSS OAI21_X1 
XU272 n157 speed[3] n1500 VDD VSS NOR2_X1 
XU271 n157 n1480 n211 N72 VDD VSS OAI21_X1 
XU270 n156 speed[2] n1490 VDD VSS NOR2_X1 
XU269 n156 N70 n210 N71 VDD VSS OAI21_X1 
XU268 speed[1] speed[0] n1480 VDD VSS NOR2_X1 
XU267 n38 n33 n39 n106 VDD VSS NAND3_X1 
XU266 state[0] n38 state[2] n730 VDD VSS NAND3_X1 
XU265 n39 n33 state[1] n700 VDD VSS NAND3_X1 
XU264 N70 n210 n211 n327 n120 VDD VSS NAND4_X1 
XU263 n213 n155 n311 n298 n119 VDD VSS NAND4_X1 
XU262 n119 n120 n118 VDD VSS NOR2_X1 
XU261 n720 n118 n730 n83 VDD VSS OAI21_X1 
XU260 n39 n38 state[2] n720 VDD VSS NAND3_X1 
XU259 state[1] state[2] n39 n64 VDD VSS NOR3_X1 
XU258 speed[6] r116_carry[6] r116_carry[7] VDD VSS OR2_X1 
XU257 speed[5] r116_carry[5] r116_carry[6] VDD VSS OR2_X1 
XU256 speed[4] r116_carry[4] r116_carry[5] VDD VSS OR2_X1 
XU255 speed[3] r116_carry[3] r116_carry[4] VDD VSS OR2_X1 
XU254 speed[2] speed[1] r116_carry[3] VDD VSS OR2_X1 
XU253 n180 n220 VDD VSS INV_X1 
XU252 n187 n221 VDD VSS INV_X1 
XSPARE_PREFIX_NAME_0 VSS VSS NETTRAN_DUMMY_2 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_1 VSS VSS NETTRAN_DUMMY_3 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_2 VSS VSS NETTRAN_DUMMY_4 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_3 VSS VSS NETTRAN_DUMMY_5 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_4 VSS VSS NETTRAN_DUMMY_6 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_5 VSS VSS NETTRAN_DUMMY_7 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_6 VSS VSS NETTRAN_DUMMY_8 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_7 VSS VSS NETTRAN_DUMMY_9 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_8 VSS VSS NETTRAN_DUMMY_10 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_9 VSS VSS NETTRAN_DUMMY_11 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_10 VSS VSS NETTRAN_DUMMY_12 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_11 VSS VSS NETTRAN_DUMMY_13 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_12 VSS VSS NETTRAN_DUMMY_14 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_13 VSS VSS NETTRAN_DUMMY_15 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_14 VSS VSS NETTRAN_DUMMY_16 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_15 VSS VSS NETTRAN_DUMMY_17 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_16 VSS VSS NETTRAN_DUMMY_18 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_17 VSS VSS NETTRAN_DUMMY_19 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_18 VSS VSS NETTRAN_DUMMY_20 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_19 VSS VSS NETTRAN_DUMMY_21 VDD VSS NOR2_X4 
XSPARE_PREFIX_NAME_0_0 VSS VSS NETTRAN_DUMMY_22 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_1 VSS VSS NETTRAN_DUMMY_23 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_2 VSS VSS NETTRAN_DUMMY_24 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_3 VSS VSS NETTRAN_DUMMY_25 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_4 VSS VSS NETTRAN_DUMMY_26 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_5 VSS VSS NETTRAN_DUMMY_27 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_6 VSS VSS NETTRAN_DUMMY_28 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_7 VSS VSS NETTRAN_DUMMY_29 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_8 VSS VSS NETTRAN_DUMMY_30 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_9 VSS VSS NETTRAN_DUMMY_31 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_10 VSS VSS NETTRAN_DUMMY_32 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_11 VSS VSS NETTRAN_DUMMY_33 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_12 VSS VSS NETTRAN_DUMMY_34 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_13 VSS VSS NETTRAN_DUMMY_35 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_14 VSS VSS NETTRAN_DUMMY_36 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_15 VSS VSS NETTRAN_DUMMY_37 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_16 VSS VSS NETTRAN_DUMMY_38 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_17 VSS VSS NETTRAN_DUMMY_39 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_18 VSS VSS NETTRAN_DUMMY_40 VDD VSS NAND2_X4 
XSPARE_PREFIX_NAME_0_19 VSS VSS NETTRAN_DUMMY_41 VDD VSS NAND2_X4 
XU114 n285 n338 VDD VSS BUF_X1 
Xadd_118 N153 N152 N151 N150 N149 N148 N147 N146 cruisespeed[7] cruisespeed[6] cruisespeed[5] 
+ cruisespeed[4] cruisespeed[3] cruisespeed[2] cruisespeed[1] cruisespeed[0] VDD 
+ VSS cruisecontrol_DW01_inc_0 
Xr113 n2 n3 n4 n5 n6 n7 n8 n9 speed[7] speed[6] speed[5] speed[4] speed[3] speed[2] 
+ speed[1] speed[0] VDD VSS cruisecontrol_DW01_inc_1 
.ENDS

